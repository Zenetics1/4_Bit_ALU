module addr (
    input wire [3:0] addr_IN,
    output wire [3:0] addr_OUT
);
    
endmodule