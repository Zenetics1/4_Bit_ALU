module subtraction(
    input wire [3:0] sub_IN,
    output wire [3:0] sub_OUT
);
    
endmodule